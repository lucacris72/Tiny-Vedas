module decode (
    input  logic        [31:0] i,
    output decode_out_t        decode_out
);
  assign decode_out.alu = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]
    &i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]&~i[12]&~i[6]&i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]
    &~i[13]&i[12]&~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&~i[12]&~i[6]&i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]
    &~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]&i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&i[2]
    &i[1]&i[0]) | (i[6]&i[5]&~i[4]&i[3]&i[2]&i[1]&i[0]) | (~i[14]&~i[13]
    &i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]
    &i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&i[12]&i[6]&i[5]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (i[14]&i[13]&i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (i[14]&i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]
    &~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[6]&~i[5]
    &i[4]&~i[3]&i[2]&i[1]&i[0]) | (~i[6]&i[5]&i[4]&~i[3]&i[2]&i[1]&i[0]) | (
    ~i[14]&i[13]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.rs1 = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&~i[5]&~i[4]&i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&~i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]&i[12]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&~i[25]&i[14]&i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]
    &~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]
    &~i[25]&i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&i[14]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&i[25]&~i[14]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]
    &~i[4]&~i[3]&i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[12]&~i[6]&~i[5]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&i[12]&i[6]&i[5]&~i[4]&~i[3]
    &~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[14]&~i[13]&i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[14]&~i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[12]
    &i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&i[13]&i[12]&~i[6]
    &~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&i[13]&~i[12]&~i[6]&~i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[12]&~i[6]&i[5]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]
    &~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]
    &i[13]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.rs2 = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&~i[5]&~i[4]&i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]
    &i[14]&i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]
    &~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]&~i[12]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]
    &~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&i[14]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&i[25]&~i[14]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&i[12]&i[6]&i[5]
    &~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&i[12]&~i[6]&i[5]&~i[4]&~i[3]
    &~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (i[14]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]
    &~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.imm12 = (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&i[2]&i[1]&i[0]) | (
    i[14]&i[13]&i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]
    &i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[13]
    &~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]
    &~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[6]
    &~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.rd = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&~i[5]&~i[4]&i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&~i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]
    &~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]&i[12]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&~i[25]&i[14]&i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[31]&i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]
    &~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]&~i[6]&i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]
    &~i[25]&i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&i[14]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]&~i[28]
    &~i[27]&~i[26]&i[25]&~i[14]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]
    &~i[4]&~i[3]&i[2]&i[1]&i[0]) | (i[6]&i[5]&~i[4]&i[3]&i[2]&i[1]&i[0]) | (
    ~i[14]&i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&i[13]&i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]
    &i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]
    &~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&i[12]&~i[6]
    &~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&~i[12]&~i[6]&~i[5]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[6]&~i[5]&i[4]&~i[3]&i[2]&i[1]&i[0]) | (~i[6]&i[5]
    &i[4]&~i[3]&i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[6]&~i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]);

  assign decode_out.shimm5 = (~i[31]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]
    &~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&~i[5]&i[4]
    &~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.imm20 = (i[6]&i[5]&~i[4]&i[3]&i[2]&i[1]&i[0]) | (~i[6]&~i[5]&i[4]&~i[3]
    &i[2]&i[1]&i[0]) | (~i[6]&i[5]&i[4]&~i[3]&i[2]&i[1]&i[0]);

  assign decode_out.pc = (i[6]&i[5]&~i[4]&i[3]&i[2]&i[1]&i[0]) | (~i[6]&~i[5]&i[4]&~i[3]&i[2]
    &i[1]&i[0]);

  assign decode_out.load = (~i[14]&i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[13]&i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&~i[12]
    &~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.store = (~i[14]&~i[13]&i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&~i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.lsu = (~i[14]&i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&~i[13]&i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]
    &~i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]
    &i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&i[12]
    &~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[13]&~i[12]&~i[6]&~i[5]
    &~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.add = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]
    &~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[6]&~i[5]&i[4]&~i[3]
    &i[2]&i[1]&i[0]);

  assign decode_out.sub = (~i[31]&i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[14]&~i[13]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]
    &i[0]) | (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    i[14]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[12]
    &i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[6]&~i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.land = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]
    &i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&i[13]&i[12]
    &~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.lor = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&i[13]&~i[12]
    &~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&i[13]&~i[12]&~i[6]
    &~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[6]&i[5]&i[4]&~i[3]&i[2]&i[1]
    &i[0]);

  assign decode_out.lxor = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]
    &~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[13]&~i[12]
    &~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.sll = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]);

  assign decode_out.sra = (~i[31]&i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]&i[12]
    &~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.srl = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&i[14]&~i[13]
    &i[12]&~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.slt = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&i[13]&~i[6]&~i[5]&i[4]
    &~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.unsign = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&i[13]
    &i[12]&~i[6]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&i[25]&i[14]&i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (i[14]&i[13]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&i[13]&i[12]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]
    &~i[13]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.condbr = (~i[14]&~i[13]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]
    &i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[14]&~i[12]&i[6]
    &i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.beq = (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.bne = (~i[14]&~i[13]&i[12]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.bge = (i[14] & i[12] & i[6] & i[5] & ~i[4] & ~i[3] & ~i[2] & i[1] & i[0]);

  assign decode_out.blt = (i[14] & ~i[12] & i[6] & i[5] & ~i[4] & ~i[3] & ~i[2] & i[1] & i[0]);

  assign decode_out.jal = (~i[14]&~i[13]&~i[12]&i[6]&i[5]&~i[4]&~i[3]&i[2]&i[1]&i[0]) | (
    i[6]&i[5]&~i[4]&i[3]&i[2]&i[1]&i[0]);

  assign decode_out.by = (~i[14]&~i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.half = (~i[14]&~i[13]&i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[13]&i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.word = (~i[14]&i[13]&~i[12]&~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (
    ~i[14]&i[13]&~i[12]&~i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.mul = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&~i[14]&~i[6]&i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.rs1_sign = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&~i[14]&i[13]
    &~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&i[25]&~i[14]&~i[13]&i[12]&~i[6]&i[5]&i[4]&~i[3]
    &~i[2]&i[1]&i[0]);

  assign decode_out.rs2_sign = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&~i[14]&~i[13]
    &i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.low = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.div = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&i[14]&~i[6]&i[5]
    &i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.rem = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&i[25]&i[14]&i[13]&~i[6]
    &i[5]&i[4]&~i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.mac = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &i[12]&~i[6]&~i[5]&~i[4]&i[3]&~i[2]&i[1]&i[0]) | (~i[31]&~i[30]&~i[29]
    &~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&~i[12]&~i[6]&~i[5]&~i[4]
    &i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.macrst = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &i[12]&~i[6]&~i[5]&~i[4]&i[3]&~i[2]&i[1]&i[0]);

  assign decode_out.nop = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[24]&~i[23]
    &~i[22]&~i[21]&~i[20]&~i[19]&~i[18]&~i[17]&~i[16]&~i[15]&~i[14]&~i[13]
    &~i[12]&~i[11]&~i[10]&~i[9]&~i[8]&~i[7]&~i[6]&~i[5]&i[4]&~i[3]&~i[2]
    &i[1]&i[0]);

  assign decode_out.legal = (~i[31]&~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[6]&i[4]&~i[3]
    &i[1]&i[0]) | (~i[31]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]
    &~i[12]&~i[6]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[13]&~i[12]&i[6]
    &i[5]&~i[4]&~i[3]&i[1]&i[0]) | (~i[14]&~i[13]&i[5]&~i[4]&~i[3]&~i[2]
    &i[1]&i[0]) | (~i[12]&~i[6]&~i[5]&i[4]&~i[3]&i[1]&i[0]) | (~i[31]
    &~i[30]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]&~i[14]&~i[13]&~i[6]&~i[5]
    &~i[4]&~i[2]&i[1]&i[0]) | (~i[31]&~i[29]&~i[28]&~i[27]&~i[26]&~i[25]
    &i[14]&~i[13]&i[12]&~i[6]&i[4]&~i[3]&i[1]&i[0]) | (~i[31]&~i[30]
    &~i[29]&~i[28]&~i[27]&~i[26]&~i[6]&i[5]&i[4]&~i[3]&i[1]&i[0]) | (
    i[14]&i[6]&i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (i[6]&i[5]&~i[4]&i[3]
    &i[2]&i[1]&i[0]) | (i[13]&~i[6]&~i[5]&i[4]&~i[3]&i[1]&i[0]) | (~i[13]
    &~i[6]&~i[5]&~i[4]&~i[3]&~i[2]&i[1]&i[0]) | (~i[14]&~i[12]&~i[6]&~i[4]
    &~i[3]&~i[2]&i[1]&i[0]) | (~i[6]&i[4]&~i[3]&i[2]&i[1]&i[0]);

endmodule
